package package_types is
  type function_select is (ADD_n, SUB_n, MUL_n, DIV_n, LSL_n, LSR_n, ASR_n, AND_n, NAND_n, NOR_n, XNOR_N, XOR_n, OR_n, ROTR_n, ROTL_n)
  
end package package_types;
 
-- Package Body
--package body package_types is
--end package body package_types;
